
module final(
    input clk;
    output reg [15:0] saida;
);

    // junção do BC com BO

    BC bc_0();

    BO bo_0();



endmodule