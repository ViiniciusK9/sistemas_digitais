
module final(output reg [15:0] saida;);



endmodule